// interface.sv

interface test_interface(input logic clk);

	// input_1
	logic	[7:0]	input_1;
	// input_2
	logic 	[7:0]	input_2;

	// output_1
	logic	[15:0]	output_1;

endinterface
